* NGSPICE file created from goldwin_dff_v2.ext - technology: sky130A

.subckt goldwin_nand_v2 A B Y VP VN
X0 Y B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
**devattr s=10000,300 d=18000,580
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=10000,300
X2 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=30000,700
X3 VP B Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
**devattr s=30000,700 d=54000,1380
.ends

.subckt goldwin_not_v2 A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=54000,1380
.ends

.subckt goldwin_dff_v2 D CLK Q QI VP VN
Xgoldwin_nand_v2_0 goldwin_nand_v2_1/Y QI Q VP VN goldwin_nand_v2
Xgoldwin_nand_v2_1 CLK D goldwin_nand_v2_1/Y VP VN goldwin_nand_v2
Xgoldwin_nand_v2_2 goldwin_nand_v2_3/Y Q QI VP VN goldwin_nand_v2
Xgoldwin_nand_v2_3 goldwin_not_v2_0/Y CLK goldwin_nand_v2_3/Y VP VN goldwin_nand_v2
Xgoldwin_not_v2_0 D goldwin_not_v2_0/Y VP VN goldwin_not_v2
.ends

