* PEX produced on Sun Apr 20 07:42:41 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_and.ext - technology: sky130A

.subckt goldwin_and A B Y VP VN
X0 a_30_540# B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X2 Y a_30_540# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
X3 a_30_540# A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X4 Y a_30_540# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
X5 VP B a_30_540# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
C0 a_30_540# a_30_0# 0.05569f
C1 B A 0.15942f
C2 Y VP 0.23897f
C3 Y a_30_540# 0.09631f
C4 B VP 0.08037f
C5 B a_30_0# 0.02784f
C6 B a_30_540# 0.13804f
C7 A VP 0.14585f
C8 A a_30_540# 0.05141f
C9 a_30_540# VP 0.53763f
C10 Y VN 0.37689f
C11 B VN 0.38251f
C12 A VN 0.37097f
C13 VP VN 2.11644f
C14 a_30_0# VN 0.0876f
C15 a_30_540# VN 0.62024f
.ends

