magic
tech sky130A
timestamp 1745127950
<< nwell >>
rect -65 250 145 645
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
<< pmos >>
rect 0 270 15 570
rect 65 270 80 570
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 125 100
rect 80 15 95 85
rect 115 15 125 85
rect 80 0 125 15
<< pdiff >>
rect -45 555 0 570
rect -45 485 -35 555
rect -15 485 0 555
rect -45 455 0 485
rect -45 385 -35 455
rect -15 385 0 455
rect -45 355 0 385
rect -45 285 -35 355
rect -15 285 0 355
rect -45 270 0 285
rect 15 555 65 570
rect 15 485 30 555
rect 50 485 65 555
rect 15 455 65 485
rect 15 385 30 455
rect 50 385 65 455
rect 15 355 65 385
rect 15 285 30 355
rect 50 285 65 355
rect 15 270 65 285
rect 80 555 125 570
rect 80 485 95 555
rect 115 485 125 555
rect 80 455 125 485
rect 80 385 95 455
rect 115 385 125 455
rect 80 355 125 385
rect 80 285 95 355
rect 115 285 125 355
rect 80 270 125 285
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
<< pdiffc >>
rect -35 485 -15 555
rect -35 385 -15 455
rect -35 285 -15 355
rect 30 485 50 555
rect 30 385 50 455
rect 30 285 50 355
rect 95 485 115 555
rect 95 385 115 455
rect 95 285 115 355
<< psubdiff >>
rect -45 -55 -25 -35
rect -5 -55 125 -35
<< nsubdiff >>
rect -45 605 -25 625
rect -5 605 85 625
rect 105 605 125 625
<< psubdiffcont >>
rect -25 -55 -5 -35
<< nsubdiffcont >>
rect -25 605 -5 625
rect 85 605 105 625
<< poly >>
rect 0 570 15 585
rect 65 570 80 585
rect 0 240 15 270
rect -5 235 15 240
rect -45 230 15 235
rect -45 210 -35 230
rect -15 210 15 230
rect -45 205 15 210
rect -5 200 15 205
rect 0 100 15 200
rect 65 165 80 270
rect 40 160 80 165
rect 40 140 50 160
rect 70 140 80 160
rect 40 135 80 140
rect 65 100 80 135
rect 0 -15 15 0
rect 65 -15 80 0
<< polycont >>
rect -35 210 -15 230
rect 50 140 70 160
<< locali >>
rect -25 625 -5 635
rect -25 560 -5 605
rect 85 625 105 635
rect 85 560 105 605
rect -45 555 -5 560
rect -45 485 -35 555
rect -15 485 -5 555
rect -45 455 -5 485
rect -45 385 -35 455
rect -15 385 -5 455
rect -45 355 -5 385
rect -45 285 -35 355
rect -15 285 -5 355
rect -45 280 -5 285
rect 20 555 60 560
rect 20 485 30 555
rect 50 485 60 555
rect 20 455 60 485
rect 20 385 30 455
rect 50 385 60 455
rect 20 355 60 385
rect 20 285 30 355
rect 50 285 60 355
rect 20 280 60 285
rect 85 555 125 560
rect 85 485 95 555
rect 115 485 125 555
rect 85 455 125 485
rect 85 385 95 455
rect 115 385 125 455
rect 85 355 125 385
rect 85 285 95 355
rect 115 285 125 355
rect 85 280 125 285
rect -45 230 -5 240
rect -45 210 -35 230
rect -15 210 -5 230
rect 30 230 50 280
rect 85 230 125 240
rect 30 210 95 230
rect 115 210 125 230
rect -45 200 -5 210
rect 85 200 125 210
rect -45 160 -5 170
rect 40 160 80 165
rect -45 140 -35 160
rect -15 140 50 160
rect 70 140 80 160
rect -45 130 -5 140
rect 40 135 80 140
rect 105 90 125 200
rect -45 85 -5 90
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect 85 85 125 90
rect 85 15 95 85
rect 115 15 125 85
rect 85 10 125 15
rect -25 -35 -5 10
rect -25 -65 -5 -55
<< viali >>
rect -25 605 -5 625
rect 85 605 105 625
rect -35 210 -15 230
rect 95 210 115 230
rect -35 140 -15 160
rect -25 -55 -5 -35
<< metal1 >>
rect -65 625 145 635
rect -65 605 -25 625
rect -5 605 85 625
rect 105 605 145 625
rect -65 595 145 605
rect -45 230 -5 240
rect -45 210 -35 230
rect -15 210 -5 230
rect -45 200 -5 210
rect 85 230 125 240
rect 85 210 95 230
rect 115 210 125 230
rect 85 200 125 210
rect -45 160 -5 170
rect -45 140 -35 160
rect -15 140 -5 160
rect -45 130 -5 140
rect -65 -35 145 -25
rect -65 -55 -25 -35
rect -5 -55 145 -35
rect -65 -65 145 -55
<< labels >>
flabel metal1 125 595 145 625 1 FreeSans 200 0 0 -120 VP
port 4 n
flabel metal1 125 -55 145 -25 1 FreeSans 200 0 0 -120 VN
port 5 n
flabel metal1 85 200 125 240 1 FreeSans 200 0 0 -120 Y
port 3 n
flabel metal1 -45 200 -5 240 1 FreeSans 200 0 0 -120 A
port 1 n
flabel metal1 -45 130 -5 170 1 FreeSans 200 0 0 -120 B
port 2 n
<< end >>
