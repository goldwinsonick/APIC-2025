* PEX produced on Sun Apr 20 09:54:23 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_dff_v2.ext - technology: sky130A

.subckt goldwin_dff_v2 D CLK Q QI VP VN
X0 goldwin_nand_v2_1.Y D a_450_n380# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X1 a_450_n380# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X2 goldwin_nand_v2_3.Y CLK a_450_120# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X3 VP CLK goldwin_nand_v2_3.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X4 goldwin_nand_v2_1.Y CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X5 a_450_120# goldwin_not_v2_0.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X6 goldwin_nand_v2_3.Y goldwin_not_v2_0.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X7 Q goldwin_nand_v2_1.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X8 VP D goldwin_nand_v2_1.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X9 Q QI a_870_n380# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X10 QI Q a_870_120# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X11 VP Q QI VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X12 VP QI Q VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X13 a_870_120# goldwin_nand_v2_3.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X14 QI goldwin_nand_v2_3.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X15 a_870_n380# goldwin_nand_v2_1.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X16 goldwin_not_v2_0.Y D VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X17 goldwin_not_v2_0.Y D VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
C0 goldwin_not_v2_0.Y goldwin_nand_v2_3.Y 0.09157f
C1 goldwin_nand_v2_1.Y Q 0.09362f
C2 QI D 0.01253f
C3 VP Q 0.63063f
C4 Q a_870_120# 0.03858f
C5 CLK goldwin_not_v2_0.Y 0.31635f
C6 a_450_n380# CLK 0.0123f
C7 CLK D 0.73431f
C8 a_870_n380# QI 0.05509f
C9 a_450_n380# goldwin_nand_v2_1.Y 0.05569f
C10 goldwin_nand_v2_1.Y D 0.14529f
C11 QI goldwin_nand_v2_3.Y 0.12351f
C12 VP goldwin_not_v2_0.Y 0.55444f
C13 VP D 0.3023f
C14 CLK goldwin_nand_v2_3.Y 0.14909f
C15 goldwin_nand_v2_3.Y a_450_120# 0.05569f
C16 a_870_n380# Q 0.05836f
C17 CLK a_450_120# 0.03278f
C18 QI goldwin_nand_v2_1.Y 0.19601f
C19 VP goldwin_nand_v2_3.Y 0.71775f
C20 VP QI 0.87457f
C21 QI a_870_120# 0.07267f
C22 goldwin_not_v2_0.Y D 0.16629f
C23 Q goldwin_nand_v2_3.Y 0.19091f
C24 goldwin_nand_v2_1.Y CLK 0.08225f
C25 a_450_n380# D 0.02784f
C26 QI Q 0.86766f
C27 VP CLK 0.38559f
C28 CLK Q 0.01253f
C29 VP goldwin_nand_v2_1.Y 0.72097f
C30 QI VN 0.7671f
C31 Q VN 0.98217f
C32 CLK VN 0.99287f
C33 D VN 1.16231f
C34 VP VN 7.49373f
C35 a_870_n380# VN 0.08205f
C36 a_450_n380# VN 0.0825f
C37 goldwin_nand_v2_1.Y VN 0.46165f
C38 a_870_120# VN 0.08205f
C39 a_450_120# VN 0.0825f
C40 goldwin_nand_v2_3.Y VN 0.44414f
C41 goldwin_not_v2_0.Y VN 0.49505f
.ends

