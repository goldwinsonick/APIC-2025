* PEX produced on Sun Apr 20 09:54:20 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_not_v2.ext - technology: sky130A

.subckt goldwin_not_v2 A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
C0 Y A 0.12139f
C1 VP A 0.12917f
C2 Y VP 0.23959f
C3 Y VN 0.39776f
C4 A VN 0.39978f
C5 VP VN 0.90177f
.ends

