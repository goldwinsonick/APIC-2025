* PEX produced on Sun Apr 20 07:42:38 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_not.ext - technology: sky130A

.subckt goldwin_not A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
C0 Y A 0.09689f
C1 VP A 0.14673f
C2 Y VP 0.23595f
C3 Y VN 0.40157f
C4 A VN 0.44806f
C5 VP VN 1.0067f
.ends

