magic
tech sky130A
timestamp 1744434067
<< nwell >>
rect -105 250 325 590
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
rect 240 0 255 100
<< pmos >>
rect 0 270 15 570
rect 65 270 80 570
rect 240 270 255 570
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 125 100
rect 80 15 95 85
rect 115 15 125 85
rect 80 0 125 15
rect 195 85 240 100
rect 195 15 205 85
rect 225 15 240 85
rect 195 0 240 15
rect 255 85 305 100
rect 255 15 270 85
rect 290 15 305 85
rect 255 0 305 15
<< pdiff >>
rect -45 555 0 570
rect -45 485 -35 555
rect -15 485 0 555
rect -45 455 0 485
rect -45 385 -35 455
rect -15 385 0 455
rect -45 355 0 385
rect -45 285 -35 355
rect -15 285 0 355
rect -45 270 0 285
rect 15 555 65 570
rect 15 485 30 555
rect 50 485 65 555
rect 15 455 65 485
rect 15 385 30 455
rect 50 385 65 455
rect 15 355 65 385
rect 15 285 30 355
rect 50 285 65 355
rect 15 270 65 285
rect 80 555 125 570
rect 80 485 95 555
rect 115 485 125 555
rect 80 455 125 485
rect 80 385 95 455
rect 115 385 125 455
rect 80 355 125 385
rect 80 285 95 355
rect 115 285 125 355
rect 80 270 125 285
rect 195 555 240 570
rect 195 485 205 555
rect 225 485 240 555
rect 195 455 240 485
rect 195 385 205 455
rect 225 385 240 455
rect 195 355 240 385
rect 195 285 205 355
rect 225 285 240 355
rect 195 270 240 285
rect 255 555 305 570
rect 255 485 270 555
rect 290 485 305 555
rect 255 455 305 485
rect 255 385 270 455
rect 290 385 305 455
rect 255 355 305 385
rect 255 285 270 355
rect 290 285 305 355
rect 255 270 305 285
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 205 15 225 85
rect 270 15 290 85
<< pdiffc >>
rect -35 485 -15 555
rect -35 385 -15 455
rect -35 285 -15 355
rect 30 485 50 555
rect 30 385 50 455
rect 30 285 50 355
rect 95 485 115 555
rect 95 385 115 455
rect 95 285 115 355
rect 205 485 225 555
rect 205 385 225 455
rect 205 285 225 355
rect 270 485 290 555
rect 270 385 290 455
rect 270 285 290 355
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
rect 155 85 195 100
rect 155 15 165 85
rect 185 15 195 85
rect 155 0 195 15
<< nsubdiff >>
rect -85 555 -45 570
rect -85 485 -75 555
rect -55 485 -45 555
rect -85 455 -45 485
rect -85 385 -75 455
rect -55 385 -45 455
rect -85 355 -45 385
rect -85 285 -75 355
rect -55 285 -45 355
rect -85 270 -45 285
rect 155 555 195 570
rect 155 485 165 555
rect 185 485 195 555
rect 155 455 195 485
rect 155 385 165 455
rect 185 385 195 455
rect 155 355 195 385
rect 155 285 165 355
rect 185 285 195 355
rect 155 270 195 285
<< psubdiffcont >>
rect -75 15 -55 85
rect 165 15 185 85
<< nsubdiffcont >>
rect -75 485 -55 555
rect -75 385 -55 455
rect -75 285 -55 355
rect 165 485 185 555
rect 165 385 185 455
rect 165 285 185 355
<< poly >>
rect 0 570 15 585
rect 65 570 80 585
rect 240 570 255 585
rect -85 230 -45 235
rect 0 230 15 270
rect -85 210 -75 230
rect -55 210 15 230
rect -85 205 -45 210
rect 0 100 15 210
rect 65 165 80 270
rect 40 160 80 165
rect 40 140 50 160
rect 70 140 80 160
rect 40 135 80 140
rect 170 160 210 165
rect 240 160 255 270
rect 170 140 180 160
rect 200 140 255 160
rect 170 135 210 140
rect 65 100 80 135
rect 240 100 255 140
rect 0 -15 15 0
rect 65 -15 80 0
rect 240 -15 255 0
<< polycont >>
rect -75 210 -55 230
rect 50 140 70 160
rect 180 140 200 160
<< locali >>
rect -65 620 -45 625
rect -65 560 -45 600
rect 85 620 105 625
rect 85 560 105 600
rect 175 620 195 625
rect 175 560 195 600
rect -85 555 -5 560
rect -85 485 -75 555
rect -55 485 -35 555
rect -15 485 -5 555
rect -85 455 -5 485
rect -85 385 -75 455
rect -55 385 -35 455
rect -15 385 -5 455
rect -85 355 -5 385
rect -85 285 -75 355
rect -55 285 -35 355
rect -15 285 -5 355
rect -85 280 -5 285
rect 20 555 60 560
rect 20 485 30 555
rect 50 485 60 555
rect 20 455 60 485
rect 20 385 30 455
rect 50 385 60 455
rect 20 355 60 385
rect 20 285 30 355
rect 50 285 60 355
rect 20 280 60 285
rect 85 555 125 560
rect 85 485 95 555
rect 115 485 125 555
rect 85 455 125 485
rect 85 385 95 455
rect 115 385 125 455
rect 85 355 125 385
rect 85 285 95 355
rect 115 285 125 355
rect 85 280 125 285
rect 155 555 235 560
rect 155 485 165 555
rect 185 485 205 555
rect 225 485 235 555
rect 155 455 235 485
rect 155 385 165 455
rect 185 385 205 455
rect 225 385 235 455
rect 155 355 235 385
rect 155 285 165 355
rect 185 285 205 355
rect 225 285 235 355
rect 155 280 235 285
rect 260 555 300 560
rect 260 485 270 555
rect 290 485 300 555
rect 260 455 300 485
rect 260 385 270 455
rect 290 385 300 455
rect 260 355 300 385
rect 260 285 270 355
rect 290 285 300 355
rect 260 280 300 285
rect -85 230 -45 240
rect -85 210 -75 230
rect -55 210 -45 230
rect 30 230 50 280
rect 270 240 290 280
rect 260 230 300 240
rect 30 210 125 230
rect -85 200 -45 210
rect -85 160 -45 170
rect 40 160 80 165
rect -85 140 -75 160
rect -55 140 50 160
rect 70 140 80 160
rect -85 130 -45 140
rect 40 135 80 140
rect 105 160 125 210
rect 260 210 270 230
rect 290 210 300 230
rect 260 200 300 210
rect 170 160 210 165
rect 105 140 180 160
rect 200 140 210 160
rect 105 90 125 140
rect 170 135 210 140
rect 270 90 290 200
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect 85 85 125 90
rect 85 15 95 85
rect 115 15 125 85
rect 85 10 125 15
rect 155 85 235 90
rect 155 15 165 85
rect 185 15 205 85
rect 225 15 235 85
rect 155 10 235 15
rect 260 85 300 90
rect 260 15 270 85
rect 290 15 300 85
rect 260 10 300 15
rect -65 -30 -45 10
rect -65 -55 -45 -50
rect 175 -30 195 10
rect 175 -55 195 -50
<< viali >>
rect -65 600 -45 620
rect 85 600 105 620
rect 175 600 195 620
rect -75 210 -55 230
rect -75 140 -55 160
rect 270 210 290 230
rect -65 -50 -45 -30
rect 175 -50 195 -30
<< metal1 >>
rect -105 620 325 625
rect -105 600 -65 620
rect -45 600 85 620
rect 105 600 175 620
rect 195 600 325 620
rect -105 595 325 600
rect -85 230 -45 240
rect -85 210 -75 230
rect -55 210 -45 230
rect -85 200 -45 210
rect 260 230 300 240
rect 260 210 270 230
rect 290 210 300 230
rect 260 200 300 210
rect -85 160 -45 170
rect -85 140 -75 160
rect -55 140 -45 160
rect -85 130 -45 140
rect -105 -30 325 -25
rect -105 -50 -65 -30
rect -45 -50 175 -30
rect 195 -50 325 -30
rect -105 -55 325 -50
<< labels >>
flabel metal1 305 -55 325 -25 1 FreeSans 200 0 0 -120 VN
port 5 n
flabel metal1 305 595 325 625 1 FreeSans 200 0 0 -120 VP
port 4 n
flabel metal1 265 200 295 240 1 FreeSans 200 0 0 -120 Y
port 3 n
flabel metal1 -85 200 -45 240 1 FreeSans 200 0 0 -120 A
port 1 n
flabel metal1 -85 130 -45 170 1 FreeSans 200 0 0 -120 B
port 2 n
<< end >>
