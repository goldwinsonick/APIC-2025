magic
tech sky130A
timestamp 1744467260
<< nwell >>
rect -60 305 1535 645
<< metal1 >>
rect -60 650 1535 680
rect 550 430 590 435
rect 550 400 555 430
rect 585 425 590 430
rect 1065 430 1105 435
rect 1065 425 1070 430
rect 585 405 1070 425
rect 585 400 590 405
rect 550 395 590 400
rect 1065 400 1070 405
rect 1100 400 1105 430
rect 1065 395 1105 400
rect 20 360 60 365
rect 20 330 25 360
rect 55 355 60 360
rect 635 360 675 365
rect 635 355 640 360
rect 55 335 640 355
rect 55 330 60 335
rect 20 325 60 330
rect 635 330 640 335
rect 670 330 675 360
rect 635 325 675 330
rect -40 285 0 295
rect 550 290 590 295
rect -40 265 20 285
rect -40 255 0 265
rect 165 265 205 285
rect 550 260 555 290
rect 585 260 590 290
rect 550 255 590 260
rect 635 290 675 295
rect 635 260 640 290
rect 670 260 675 290
rect 635 255 675 260
rect 980 290 1020 295
rect 980 260 985 290
rect 1015 260 1020 290
rect 980 255 1020 260
rect 1065 290 1105 295
rect 1065 260 1070 290
rect 1100 260 1105 290
rect 1475 285 1515 295
rect 1450 265 1515 285
rect 1065 255 1105 260
rect 1475 255 1515 265
rect -40 215 0 225
rect 980 220 1020 225
rect -40 195 205 215
rect -40 185 0 195
rect 980 190 985 220
rect 1015 215 1020 220
rect 1015 195 1065 215
rect 1015 190 1020 195
rect 980 185 1020 190
rect -40 145 0 155
rect 635 150 675 155
rect 635 145 640 150
rect -40 125 640 145
rect -40 115 0 125
rect 635 120 640 125
rect 670 120 675 150
rect 635 115 675 120
rect -60 0 1535 30
<< via1 >>
rect 555 400 585 430
rect 1070 400 1100 430
rect 25 330 55 360
rect 640 330 670 360
rect 25 260 55 290
rect 555 260 585 290
rect 640 260 670 290
rect 985 260 1015 290
rect 1070 260 1100 290
rect 640 190 670 220
rect 985 190 1015 220
rect 640 120 670 150
<< metal2 >>
rect 550 430 590 435
rect 550 400 555 430
rect 585 400 590 430
rect 550 395 590 400
rect 1065 430 1105 435
rect 1065 400 1070 430
rect 1100 400 1105 430
rect 1065 395 1105 400
rect 20 360 60 365
rect 20 330 25 360
rect 55 330 60 360
rect 20 325 60 330
rect 30 295 50 325
rect 560 295 580 395
rect 635 360 675 365
rect 635 330 640 360
rect 670 330 675 360
rect 635 325 675 330
rect 645 295 665 325
rect 1075 295 1095 395
rect 20 290 60 295
rect 20 260 25 290
rect 55 260 60 290
rect 20 255 60 260
rect 550 290 590 295
rect 550 260 555 290
rect 585 260 590 290
rect 550 255 590 260
rect 635 290 675 295
rect 635 260 640 290
rect 670 260 675 290
rect 635 255 675 260
rect 980 290 1020 295
rect 980 260 985 290
rect 1015 260 1020 290
rect 980 255 1020 260
rect 1065 290 1105 295
rect 1065 260 1070 290
rect 1100 260 1105 290
rect 1065 255 1105 260
rect 990 225 1010 255
rect 635 220 675 225
rect 635 190 640 220
rect 670 190 675 220
rect 635 185 675 190
rect 980 220 1020 225
rect 980 190 985 220
rect 1015 190 1020 220
rect 980 185 1020 190
rect 645 155 665 185
rect 635 150 675 155
rect 635 120 640 150
rect 670 120 675 150
rect 635 115 675 120
use goldwin_and  goldwin_and_1 ../goldwin_and
timestamp 1744434067
transform 1 0 290 0 1 55
box -105 -55 325 625
use goldwin_and  goldwin_and_2
timestamp 1744434067
transform 1 0 720 0 1 55
box -105 -55 325 625
use goldwin_not  goldwin_not_0 ../goldwin_not
timestamp 1744448201
transform 1 0 105 0 1 55
box -105 -55 80 625
use goldwin_or  goldwin_or_0 ../goldwin_or
timestamp 1744434135
transform 1 0 1150 0 1 55
box -105 -55 325 625
<< labels >>
flabel metal1 -40 185 0 225 1 FreeSans 200 0 0 -120 A
port 1 n
flabel metal1 -40 115 0 155 1 FreeSans 200 0 0 -120 B
port 2 n
flabel metal1 1475 255 1515 295 1 FreeSans 200 0 0 -120 Y
port 4 n
flabel metal1 1495 0 1515 30 1 FreeSans 200 0 0 -120 VN
port 6 n
flabel metal1 1495 650 1515 680 1 FreeSans 200 0 0 -120 VP
port 5 n
flabel metal1 -40 255 0 295 1 FreeSans 200 0 0 -120 S
port 3 n
<< end >>
