magic
tech sky130A
timestamp 1744179846
<< nwell >>
rect -80 -10 355 140
<< nmos >>
rect -10 -275 5 -175
rect 120 -275 135 -175
rect 270 -275 285 -175
<< pmos >>
rect -10 15 5 115
rect 120 15 135 115
rect 270 15 285 115
<< ndiff >>
rect -60 -245 -10 -175
rect -60 -265 -55 -245
rect -35 -265 -10 -245
rect -60 -275 -10 -265
rect 5 -185 120 -175
rect 5 -205 30 -185
rect 50 -205 120 -185
rect 5 -275 120 -205
rect 135 -185 190 -175
rect 135 -205 165 -185
rect 185 -205 190 -185
rect 135 -275 190 -205
rect 220 -245 270 -175
rect 220 -265 225 -245
rect 245 -265 270 -245
rect 220 -275 270 -265
rect 285 -185 335 -175
rect 285 -205 310 -185
rect 330 -205 335 -185
rect 285 -275 335 -205
<< pdiff >>
rect -60 105 -10 115
rect -60 85 -55 105
rect -35 85 -10 105
rect -60 15 -10 85
rect 5 45 120 115
rect 5 25 30 45
rect 50 25 120 45
rect 5 15 120 25
rect 135 110 160 115
rect 135 100 190 110
rect 135 80 165 100
rect 185 80 190 100
rect 135 15 190 80
rect 220 100 270 115
rect 220 80 225 100
rect 245 80 270 100
rect 220 15 270 80
rect 285 50 335 115
rect 285 30 310 50
rect 330 30 335 50
rect 285 15 335 30
<< ndiffc >>
rect -55 -265 -35 -245
rect 30 -205 50 -185
rect 165 -205 185 -185
rect 225 -265 245 -245
rect 310 -205 330 -185
<< pdiffc >>
rect -55 85 -35 105
rect 30 25 50 45
rect 165 80 185 100
rect 225 80 245 100
rect 310 30 330 50
<< poly >>
rect -10 115 5 140
rect 120 115 135 140
rect 270 115 285 140
rect -10 -30 5 15
rect 120 -30 135 15
rect -35 -35 5 -30
rect -35 -55 -25 -35
rect -5 -55 5 -35
rect -35 -60 5 -55
rect 95 -35 135 -30
rect 95 -55 105 -35
rect 125 -55 135 -35
rect 95 -60 135 -55
rect -10 -175 5 -60
rect 120 -175 135 -60
rect 270 -115 285 15
rect 245 -120 285 -115
rect 245 -140 255 -120
rect 275 -140 285 -120
rect 245 -145 285 -140
rect 270 -175 285 -145
rect -10 -295 5 -275
rect 120 -295 135 -275
rect 270 -295 285 -275
<< polycont >>
rect -25 -55 -5 -35
rect 105 -55 125 -35
rect 255 -140 275 -120
<< locali >>
rect -60 105 -30 115
rect -60 85 -55 105
rect -35 85 -30 105
rect -60 75 -30 85
rect 160 100 190 110
rect 160 80 165 100
rect 185 80 190 100
rect 160 70 190 80
rect 220 100 250 110
rect 220 80 225 100
rect 245 80 250 100
rect 220 70 250 80
rect 25 45 55 55
rect 25 25 30 45
rect 50 25 55 45
rect 25 15 55 25
rect 305 50 335 60
rect 305 30 310 50
rect 330 30 335 50
rect 305 20 335 30
rect -35 -35 5 -30
rect -35 -55 -25 -35
rect -5 -55 5 -35
rect -35 -60 5 -55
rect 95 -35 135 -30
rect 95 -55 105 -35
rect 125 -55 135 -35
rect 95 -60 135 -55
rect 245 -120 285 -115
rect 245 -140 255 -120
rect 275 -140 285 -120
rect 245 -145 285 -140
rect 25 -185 55 -175
rect 25 -205 30 -185
rect 50 -205 55 -185
rect 25 -215 55 -205
rect 160 -185 190 -175
rect 160 -205 165 -185
rect 185 -205 190 -185
rect 160 -215 190 -205
rect 305 -185 335 -175
rect 305 -205 310 -185
rect 330 -205 335 -185
rect 305 -215 335 -205
rect -60 -245 -30 -235
rect -60 -265 -55 -245
rect -35 -265 -30 -245
rect -60 -275 -30 -265
rect 220 -245 250 -235
rect 220 -265 225 -245
rect 245 -265 250 -245
rect 220 -275 250 -265
<< metal1 >>
rect -80 155 355 185
rect -60 85 -30 155
rect 160 80 190 155
rect 220 80 250 155
rect -55 -60 5 -30
rect 25 -115 55 55
rect 75 -60 135 -30
rect 25 -145 285 -115
rect 25 -215 55 -145
rect 160 -215 190 -145
rect 305 -215 335 60
rect -60 -310 -30 -235
rect 220 -310 250 -235
rect -80 -340 355 -310
<< end >>
