* PEX produced on Fri Apr 18 07:54:14 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_nand.ext - technology: sky130A

.subckt goldwin_nand A B Y VP VN
X0 Y B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X2 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X3 VP B Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
C0 B VP 0.07599f
C1 Y A 0.06452f
C2 B A 0.15942f
C3 Y B 0.11686f
C4 Y a_30_0# 0.05569f
C5 A VP 0.14585f
C6 Y VP 0.45643f
C7 a_30_0# B 0.02784f
C8 Y VN 0.25248f
C9 B VN 0.4103f
C10 A VN 0.36737f
C11 VP VN 1.39457f
C12 a_30_0# VN 0.08711f
.ends

