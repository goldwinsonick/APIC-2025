magic
tech sky130A
timestamp 1744474457
<< nwell >>
rect -60 305 1245 645
<< metal1 >>
rect -60 650 1245 680
rect 705 435 745 440
rect 705 405 710 435
rect 740 430 745 435
rect 1125 435 1165 440
rect 1125 430 1130 435
rect 740 410 1130 430
rect 740 405 745 410
rect 705 400 745 405
rect 1125 405 1130 410
rect 1160 405 1165 435
rect 1125 400 1165 405
rect 20 360 60 365
rect 20 330 25 360
rect 55 355 60 360
rect 455 360 495 365
rect 455 355 460 360
rect 55 335 460 355
rect 55 330 60 335
rect 20 325 60 330
rect 455 330 460 335
rect 490 330 495 360
rect 455 325 495 330
rect 625 360 665 365
rect 625 330 630 360
rect 660 355 665 360
rect 875 355 915 365
rect 955 360 995 365
rect 955 355 960 360
rect 660 335 960 355
rect 660 330 665 335
rect 625 325 665 330
rect 875 325 915 335
rect 955 330 960 335
rect 990 330 995 360
rect 955 325 995 330
rect -40 285 0 295
rect 455 290 495 295
rect -40 265 20 285
rect -40 255 0 265
rect 165 265 205 285
rect 455 260 460 290
rect 490 260 495 290
rect 455 255 495 260
rect 625 290 665 295
rect 625 260 630 290
rect 660 260 665 290
rect 625 255 665 260
rect 705 290 745 295
rect 705 260 710 290
rect 740 260 745 290
rect 705 255 745 260
rect 875 290 915 295
rect 875 260 880 290
rect 910 260 915 290
rect 875 255 915 260
rect 955 290 995 295
rect 955 260 960 290
rect 990 260 995 290
rect 955 255 995 260
rect 1125 290 1165 295
rect 1125 260 1130 290
rect 1160 285 1165 290
rect 1185 285 1225 295
rect 1160 265 1225 285
rect 1160 260 1165 265
rect 1125 255 1165 260
rect 1185 255 1225 265
rect -40 215 0 225
rect 875 220 915 225
rect -40 195 205 215
rect 245 195 455 215
rect -40 185 0 195
rect 875 190 880 220
rect 910 215 915 220
rect 955 215 995 225
rect 1185 215 1225 225
rect 910 195 1225 215
rect 910 190 915 195
rect 875 185 915 190
rect 955 185 995 195
rect 1185 185 1225 195
rect 375 150 415 155
rect 375 120 380 150
rect 410 145 415 150
rect 705 150 745 155
rect 705 145 710 150
rect 410 125 710 145
rect 410 120 415 125
rect 375 115 415 120
rect 705 120 710 125
rect 740 120 745 150
rect 705 115 745 120
rect -60 0 1245 30
<< via1 >>
rect 710 405 740 435
rect 1130 405 1160 435
rect 25 330 55 360
rect 460 330 490 360
rect 630 330 660 360
rect 960 330 990 360
rect 25 260 55 290
rect 380 260 410 290
rect 460 260 490 290
rect 630 260 660 290
rect 710 260 740 290
rect 880 260 910 290
rect 960 260 990 290
rect 1130 260 1160 290
rect 710 190 740 220
rect 880 190 910 220
rect 380 120 410 150
rect 710 120 740 150
<< metal2 >>
rect 705 435 745 440
rect 705 405 710 435
rect 740 405 745 435
rect 705 400 745 405
rect 1125 435 1165 440
rect 1125 405 1130 435
rect 1160 405 1165 435
rect 1125 400 1165 405
rect 20 360 60 365
rect 20 330 25 360
rect 55 330 60 360
rect 20 325 60 330
rect 455 360 495 365
rect 455 330 460 360
rect 490 330 495 360
rect 455 325 495 330
rect 625 360 665 365
rect 625 330 630 360
rect 660 330 665 360
rect 625 325 665 330
rect 30 295 50 325
rect 465 295 485 325
rect 635 295 655 325
rect 715 295 735 400
rect 955 360 995 365
rect 955 330 960 360
rect 990 330 995 360
rect 955 325 995 330
rect 965 295 985 325
rect 1135 295 1155 400
rect 20 290 60 295
rect 20 260 25 290
rect 55 260 60 290
rect 20 255 60 260
rect 375 290 415 295
rect 375 260 380 290
rect 410 260 415 290
rect 375 255 415 260
rect 455 290 495 295
rect 455 260 460 290
rect 490 260 495 290
rect 455 255 495 260
rect 625 290 665 295
rect 625 260 630 290
rect 660 260 665 290
rect 625 255 665 260
rect 705 290 745 295
rect 705 260 710 290
rect 740 260 745 290
rect 705 255 745 260
rect 875 290 915 295
rect 875 260 880 290
rect 910 260 915 290
rect 875 255 915 260
rect 955 290 995 295
rect 955 260 960 290
rect 990 260 995 290
rect 955 255 995 260
rect 1125 290 1165 295
rect 1125 260 1130 290
rect 1160 260 1165 290
rect 1125 255 1165 260
rect 385 155 405 255
rect 885 225 905 255
rect 705 220 745 225
rect 705 190 710 220
rect 740 190 745 220
rect 705 185 745 190
rect 875 220 915 225
rect 875 190 880 220
rect 910 190 915 220
rect 875 185 915 190
rect 715 155 735 185
rect 375 150 415 155
rect 375 120 380 150
rect 410 120 415 150
rect 375 115 415 120
rect 705 150 745 155
rect 705 120 710 150
rect 740 120 745 150
rect 705 115 745 120
use goldwin_nand  goldwin_nand_0 ../goldwin_nand
timestamp 1744432086
transform 1 0 1040 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_1
timestamp 1744432086
transform 1 0 290 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_2
timestamp 1744432086
transform 1 0 540 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_3
timestamp 1744432086
transform 1 0 790 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_4
timestamp 1744432086
transform 1 0 790 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_5
timestamp 1744432086
transform 1 0 540 0 1 55
box -105 -55 145 625
use goldwin_nand  goldwin_nand_6
timestamp 1744432086
transform 1 0 290 0 1 55
box -105 -55 145 625
use goldwin_not  goldwin_not_0 ../goldwin_not
timestamp 1744448201
transform 1 0 105 0 1 55
box -105 -55 80 625
<< labels >>
flabel metal1 -40 255 0 295 1 FreeSans 200 0 0 -120 D
port 1 n
flabel metal1 -40 185 0 225 1 FreeSans 200 0 0 -120 CLK
port 2 n
flabel metal1 1185 255 1225 295 1 FreeSans 200 0 0 -120 Q
port 3 n
flabel metal1 1185 185 1225 225 1 FreeSans 200 0 0 -120 QI
port 4 n
flabel metal1 1205 650 1225 680 1 FreeSans 200 0 0 -120 VP
port 5 n
flabel metal1 1205 0 1225 30 1 FreeSans 200 0 0 -120 VN
port 6 n
<< end >>
