magic
tech sky130A
timestamp 1744219405
<< nwell >>
rect -120 205 305 560
<< nmos >>
rect -15 0 0 100
rect 50 0 65 100
rect 225 0 240 100
<< pmos >>
rect -15 225 0 540
rect 50 225 65 540
rect 225 225 240 540
<< ndiff >>
rect -60 85 -15 100
rect -60 15 -50 85
rect -30 15 -15 85
rect -60 0 -15 15
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 85 110 100
rect 65 15 80 85
rect 100 15 110 85
rect 65 0 110 15
rect 180 85 225 100
rect 180 15 190 85
rect 210 15 225 85
rect 180 0 225 15
rect 240 85 285 100
rect 240 15 255 85
rect 275 15 285 85
rect 240 0 285 15
<< pdiff >>
rect -60 525 -15 540
rect -60 450 -50 525
rect -30 450 -15 525
rect -60 420 -15 450
rect -60 345 -50 420
rect -30 345 -15 420
rect -60 315 -15 345
rect -60 240 -50 315
rect -30 240 -15 315
rect -60 225 -15 240
rect 0 525 50 540
rect 0 450 15 525
rect 35 450 50 525
rect 0 420 50 450
rect 0 345 15 420
rect 35 345 50 420
rect 0 315 50 345
rect 0 240 15 315
rect 35 240 50 315
rect 0 225 50 240
rect 65 525 110 540
rect 65 450 80 525
rect 100 450 110 525
rect 65 420 110 450
rect 65 345 80 420
rect 100 345 110 420
rect 65 315 110 345
rect 65 240 80 315
rect 100 240 110 315
rect 65 225 110 240
rect 180 525 225 540
rect 180 450 190 525
rect 210 450 225 525
rect 180 420 225 450
rect 180 345 190 420
rect 210 345 225 420
rect 180 315 225 345
rect 180 240 190 315
rect 210 240 225 315
rect 180 225 225 240
rect 240 525 285 540
rect 240 450 255 525
rect 275 450 285 525
rect 240 420 285 450
rect 240 345 255 420
rect 275 345 285 420
rect 240 315 285 345
rect 240 240 255 315
rect 275 240 285 315
rect 240 225 285 240
<< ndiffc >>
rect -50 15 -30 85
rect 15 15 35 85
rect 80 15 100 85
rect 190 15 210 85
rect 255 15 275 85
<< pdiffc >>
rect -50 450 -30 525
rect -50 345 -30 420
rect -50 240 -30 315
rect 15 450 35 525
rect 15 345 35 420
rect 15 240 35 315
rect 80 450 100 525
rect 80 345 100 420
rect 80 240 100 315
rect 190 450 210 525
rect 190 345 210 420
rect 190 240 210 315
rect 255 450 275 525
rect 255 345 275 420
rect 255 240 275 315
<< psubdiff >>
rect -100 85 -60 100
rect -100 15 -90 85
rect -70 15 -60 85
rect -100 0 -60 15
rect 140 85 180 100
rect 140 15 150 85
rect 170 15 180 85
rect 140 0 180 15
<< nsubdiff >>
rect -100 525 -60 540
rect -100 450 -90 525
rect -70 450 -60 525
rect -100 420 -60 450
rect -100 345 -90 420
rect -70 345 -60 420
rect -100 315 -60 345
rect -100 240 -90 315
rect -70 240 -60 315
rect -100 225 -60 240
rect 140 525 180 540
rect 140 450 150 525
rect 170 450 180 525
rect 140 420 180 450
rect 140 345 150 420
rect 170 345 180 420
rect 140 315 180 345
rect 140 240 150 315
rect 170 240 180 315
rect 140 225 180 240
<< psubdiffcont >>
rect -90 15 -70 85
rect 150 15 170 85
<< nsubdiffcont >>
rect -90 450 -70 525
rect -90 345 -70 420
rect -90 240 -70 315
rect 150 450 170 525
rect 150 345 170 420
rect 150 240 170 315
<< poly >>
rect -15 540 0 555
rect 50 540 65 555
rect 225 540 240 555
rect -15 190 0 225
rect -55 185 0 190
rect -55 165 -45 185
rect -25 165 0 185
rect -55 160 0 165
rect -15 100 0 160
rect 50 190 65 225
rect 50 185 105 190
rect 50 165 75 185
rect 95 165 105 185
rect 50 160 105 165
rect 50 100 65 160
rect 225 150 240 225
rect 185 145 240 150
rect 185 125 195 145
rect 215 125 240 145
rect 185 120 240 125
rect 225 100 240 120
rect -15 -15 0 0
rect 50 -15 65 0
rect 225 -15 240 0
<< polycont >>
rect -45 165 -25 185
rect 75 165 95 185
rect 195 125 215 145
<< locali >>
rect -100 565 -80 570
rect -100 530 -80 545
rect 90 565 110 570
rect 90 530 110 545
rect -100 525 -20 530
rect -100 450 -90 525
rect -70 450 -50 525
rect -30 450 -20 525
rect -100 445 -20 450
rect 5 525 45 530
rect 5 450 15 525
rect 35 450 45 525
rect 5 445 45 450
rect 70 525 110 530
rect 70 450 80 525
rect 100 450 110 525
rect 70 445 110 450
rect 140 565 160 570
rect 140 530 160 545
rect 140 525 220 530
rect 140 450 150 525
rect 170 450 190 525
rect 210 450 220 525
rect 140 445 220 450
rect 245 525 285 530
rect 245 450 255 525
rect 275 450 285 525
rect 245 445 285 450
rect -100 420 -20 425
rect -100 345 -90 420
rect -70 345 -50 420
rect -30 345 -20 420
rect -100 340 -20 345
rect 5 420 45 425
rect 5 345 15 420
rect 35 345 45 420
rect 5 340 45 345
rect 70 420 110 425
rect 70 345 80 420
rect 100 345 110 420
rect 70 340 110 345
rect 140 420 220 425
rect 140 345 150 420
rect 170 345 190 420
rect 210 345 220 420
rect 140 340 220 345
rect 245 420 285 425
rect 245 345 255 420
rect 275 345 285 420
rect 245 340 285 345
rect -100 315 -20 320
rect -100 240 -90 315
rect -70 240 -50 315
rect -30 240 -20 315
rect -100 235 -20 240
rect 5 315 45 320
rect 5 240 15 315
rect 35 240 45 315
rect 5 235 45 240
rect 70 315 110 320
rect 70 240 80 315
rect 100 240 110 315
rect 70 235 110 240
rect 140 315 220 320
rect 140 240 150 315
rect 170 240 190 315
rect 210 240 220 315
rect 140 235 220 240
rect 245 315 285 320
rect 245 240 255 315
rect 275 240 285 315
rect 245 235 285 240
rect -55 185 -15 190
rect -55 165 -45 185
rect -25 165 -15 185
rect -55 160 -15 165
rect 15 140 35 235
rect 255 190 275 235
rect 65 185 105 190
rect 65 165 75 185
rect 95 165 105 185
rect 65 160 105 165
rect 255 185 305 190
rect 255 165 275 185
rect 295 165 305 185
rect 255 160 305 165
rect 185 145 225 150
rect 185 140 195 145
rect 15 125 195 140
rect 215 125 225 145
rect 15 120 225 125
rect 15 90 35 120
rect 80 90 100 120
rect 255 90 275 160
rect -100 85 -20 90
rect -100 15 -90 85
rect -70 15 -50 85
rect -30 15 -20 85
rect -100 10 -20 15
rect 5 85 45 90
rect 5 15 15 85
rect 35 15 45 85
rect 5 10 45 15
rect 70 85 110 90
rect 70 15 80 85
rect 100 15 110 85
rect 70 10 110 15
rect 140 85 220 90
rect 140 15 150 85
rect 170 15 190 85
rect 210 15 220 85
rect 140 10 220 15
rect 245 85 285 90
rect 245 15 255 85
rect 275 15 285 85
rect 245 10 285 15
rect -100 -5 -80 10
rect -100 -30 -80 -25
rect 140 -5 160 10
rect 140 -30 160 -25
<< viali >>
rect -100 545 -80 565
rect 90 545 110 565
rect 140 545 160 565
rect -45 165 -25 185
rect 75 165 95 185
rect 275 165 295 185
rect -100 -25 -80 -5
rect 140 -25 160 -5
<< metal1 >>
rect -120 565 305 570
rect -120 545 -100 565
rect -80 545 90 565
rect 110 545 140 565
rect 160 545 305 565
rect -120 540 305 545
rect -120 185 -15 190
rect -120 165 -45 185
rect -25 165 -15 185
rect -120 160 -15 165
rect 65 185 145 190
rect 65 165 75 185
rect 95 165 145 185
rect 65 160 145 165
rect 255 185 305 190
rect 255 165 275 185
rect 295 165 305 185
rect 255 160 305 165
rect -120 -5 305 0
rect -120 -25 -100 -5
rect -80 -25 140 -5
rect 160 -25 305 -5
rect -120 -30 305 -25
<< labels >>
rlabel metal1 -120 175 -120 175 7 A
port 1 w
rlabel metal1 145 175 145 175 7 B
port 2 w
rlabel metal1 305 175 305 175 7 OUT
port 3 w
rlabel metal1 305 555 305 555 7 VP
port 4 w
rlabel metal1 305 -15 305 -15 7 VN
port 5 w
<< end >>
