magic
tech sky130A
timestamp 1745136940
<< nwell >>
rect -60 1045 0 1440
rect 1225 1045 1285 1440
rect -60 0 0 395
rect 1225 0 1285 395
<< metal1 >>
rect -60 1390 0 1430
rect 1225 1390 1285 1430
rect -40 1025 0 1035
rect 480 1030 520 1035
rect -40 1005 20 1025
rect -40 995 0 1005
rect 480 1000 485 1030
rect 515 1025 520 1030
rect 1225 1025 1265 1035
rect 515 1005 560 1025
rect 1205 1005 1265 1025
rect 515 1000 520 1005
rect 480 995 520 1000
rect 1225 995 1265 1005
rect -40 955 0 965
rect -40 935 20 955
rect -40 925 0 935
rect 1225 955 1265 965
rect 1205 935 1265 955
rect 1225 925 1265 935
rect -40 885 0 895
rect 560 890 600 895
rect 560 885 565 890
rect -40 865 565 885
rect -40 855 0 865
rect 560 860 565 865
rect 595 860 600 890
rect 560 855 600 860
rect -60 730 0 770
rect 1225 730 1285 770
rect -60 670 0 710
rect 1225 670 1285 710
rect 480 580 520 585
rect 480 550 485 580
rect 515 575 520 580
rect 1225 575 1265 585
rect 515 555 1265 575
rect 515 550 520 555
rect 480 545 520 550
rect 1225 545 1265 555
rect -40 435 0 445
rect 480 440 520 445
rect -40 415 20 435
rect -40 405 0 415
rect 480 410 485 440
rect 515 410 520 440
rect 480 405 520 410
rect -60 10 0 50
rect 1225 10 1285 50
<< via1 >>
rect 485 1000 515 1030
rect 565 930 595 960
rect 565 860 595 890
rect 485 550 515 580
rect 485 410 515 440
<< metal2 >>
rect 480 1030 520 1035
rect 480 1000 485 1030
rect 515 1000 520 1030
rect 480 995 520 1000
rect 490 585 510 995
rect 560 960 600 965
rect 560 930 565 960
rect 595 930 600 960
rect 560 925 600 930
rect 570 895 590 925
rect 560 890 600 895
rect 560 860 565 890
rect 595 860 600 890
rect 560 855 600 860
rect 480 580 520 585
rect 480 550 485 580
rect 515 550 520 580
rect 480 545 520 550
rect 490 445 510 545
rect 480 440 520 445
rect 480 410 485 440
rect 515 410 520 440
rect 480 405 520 410
use goldwin_dff_v2  goldwin_dff_v2_0 ../goldwin_dff_v2
timestamp 1745135597
transform 1 0 600 0 1 735
box -60 -735 625 705
use goldwin_mux_v2  goldwin_mux_v2_0 ../goldwin_mux_v2
timestamp 1745132050
transform 1 0 60 0 1 730
box -60 -730 485 710
<< labels >>
flabel metal1 -40 995 0 1035 1 FreeSans 200 0 0 0 S
port 4 n
flabel metal1 -40 925 0 965 1 FreeSans 200 0 0 0 A
port 2 n
flabel metal1 -40 855 0 895 1 FreeSans 200 0 0 0 CLK
port 1 n
flabel metal1 -40 405 0 445 1 FreeSans 200 0 0 0 B
port 3 n
flabel metal1 1225 925 1265 965 1 FreeSans 200 0 0 0 Q
port 6 n
flabel metal1 1265 1390 1285 1430 1 FreeSans 200 0 0 0 VP
port 8 n
flabel metal1 1265 730 1285 770 1 FreeSans 200 0 0 0 VN
port 9 n
flabel metal1 1225 995 1265 1035 1 FreeSans 200 0 0 0 QI
port 7 n
flabel metal1 1225 545 1265 585 1 FreeSans 200 0 0 0 D
port 5 n
<< end >>
