* NGSPICE file created from goldwin_mux_dff.ext - technology: sky130A

.subckt goldwin_and A B Y VP VN
X0 a_30_540# B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
**devattr s=10000,300 d=18000,580
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=10000,300
X2 Y a_30_540# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=20000,600
X3 a_30_540# A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=30000,700
X4 Y a_30_540# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=60000,1400
X5 VP B a_30_540# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
**devattr s=30000,700 d=54000,1380
.ends

.subckt goldwin_or A B Y VP VN
X0 VN A a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
**devattr s=10000,300 d=18000,580
X1 a_30_0# B VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=10000,300
X2 Y a_30_0# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=20000,600
X3 a_30_540# B VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=30000,700
X4 Y a_30_0# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=60000,1400
X5 a_30_0# A a_30_540# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
**devattr s=30000,700 d=54000,1380
.ends

.subckt goldwin_not A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=18000,580
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=54000,1380
.ends

.subckt goldwin_mux A B S Y VP VN
Xgoldwin_and_1 goldwin_not_0/Y A goldwin_or_0/A VP VN goldwin_and
Xgoldwin_and_2 S B goldwin_or_0/B VP VN goldwin_and
Xgoldwin_or_0 goldwin_or_0/A goldwin_or_0/B Y VP VN goldwin_or
Xgoldwin_not_0 S goldwin_not_0/Y VP VN goldwin_not
.ends

.subckt goldwin_nand A B Y VP VN a_30_0#
X0 Y B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
**devattr s=10000,300 d=18000,580
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=10000,300
X2 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
**devattr s=54000,1380 d=30000,700
X3 VP B Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
**devattr s=30000,700 d=54000,1380
.ends

.subckt goldwin_dff D CLK Q QI VP VN
Xgoldwin_nand_0 goldwin_nand_5/Y QI Q VP VN goldwin_nand_0/a_30_0# goldwin_nand
Xgoldwin_nand_1 goldwin_not_0/Y CLK goldwin_nand_6/Y VP VN goldwin_nand_6/a_30_0#
+ goldwin_nand
Xgoldwin_nand_2 D CLK goldwin_nand_5/Y VP VN goldwin_nand_5/a_30_0# goldwin_nand
Xgoldwin_nand_3 Q goldwin_nand_6/Y QI VP VN goldwin_nand_4/a_30_0# goldwin_nand
Xgoldwin_nand_4 Q goldwin_nand_6/Y QI VP VN goldwin_nand_4/a_30_0# goldwin_nand
Xgoldwin_nand_5 D CLK goldwin_nand_5/Y VP VN goldwin_nand_5/a_30_0# goldwin_nand
Xgoldwin_nand_6 goldwin_not_0/Y CLK goldwin_nand_6/Y VP VN goldwin_nand_6/a_30_0#
+ goldwin_nand
Xgoldwin_not_0 D goldwin_not_0/Y VP VN goldwin_not
.ends

.subckt goldwin_mux_dff CLK A B S D Q QI VP VN
Xgoldwin_mux_0 A B S D VP VN goldwin_mux
Xgoldwin_dff_0 D CLK Q QI VP VN goldwin_dff
.ends

