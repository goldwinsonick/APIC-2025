magic
tech sky130A
timestamp 1744448201
<< nwell >>
rect -105 250 80 590
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 270 15 570
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 60 100
rect 15 15 30 85
rect 50 15 60 85
rect 15 0 60 15
<< pdiff >>
rect -45 555 0 570
rect -45 485 -35 555
rect -15 485 0 555
rect -45 455 0 485
rect -45 385 -35 455
rect -15 385 0 455
rect -45 355 0 385
rect -45 285 -35 355
rect -15 285 0 355
rect -45 270 0 285
rect 15 555 60 570
rect 15 485 30 555
rect 50 485 60 555
rect 15 455 60 485
rect 15 385 30 455
rect 50 385 60 455
rect 15 355 60 385
rect 15 285 30 355
rect 50 285 60 355
rect 15 270 60 285
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< pdiffc >>
rect -35 485 -15 555
rect -35 385 -15 455
rect -35 285 -15 355
rect 30 485 50 555
rect 30 385 50 455
rect 30 285 50 355
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
<< nsubdiff >>
rect -85 555 -45 570
rect -85 485 -75 555
rect -55 485 -45 555
rect -85 455 -45 485
rect -85 385 -75 455
rect -55 385 -45 455
rect -85 355 -45 385
rect -85 285 -75 355
rect -55 285 -45 355
rect -85 270 -45 285
<< psubdiffcont >>
rect -75 15 -55 85
<< nsubdiffcont >>
rect -75 485 -55 555
rect -75 385 -55 455
rect -75 285 -55 355
<< poly >>
rect 0 570 15 585
rect -85 230 -45 235
rect 0 230 15 270
rect -85 210 -75 230
rect -55 210 15 230
rect -85 205 -45 210
rect 0 100 15 210
rect 0 -15 15 0
<< polycont >>
rect -75 210 -55 230
<< locali >>
rect -65 620 -45 625
rect -65 560 -45 600
rect -85 555 -5 560
rect -85 485 -75 555
rect -55 485 -35 555
rect -15 485 -5 555
rect -85 455 -5 485
rect -85 385 -75 455
rect -55 385 -35 455
rect -15 385 -5 455
rect -85 355 -5 385
rect -85 285 -75 355
rect -55 285 -35 355
rect -15 285 -5 355
rect -85 280 -5 285
rect 20 555 60 560
rect 20 485 30 555
rect 50 485 60 555
rect 20 455 60 485
rect 20 385 30 455
rect 50 385 60 455
rect 20 355 60 385
rect 20 285 30 355
rect 50 285 60 355
rect 20 280 60 285
rect 30 240 50 280
rect -85 230 -45 240
rect -85 210 -75 230
rect -55 210 -45 230
rect -85 200 -45 210
rect 20 230 60 240
rect 20 210 30 230
rect 50 210 60 230
rect 20 200 60 210
rect 30 90 50 200
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect -65 -30 -45 10
rect -65 -55 -45 -50
<< viali >>
rect -65 600 -45 620
rect -75 210 -55 230
rect 30 210 50 230
rect -65 -50 -45 -30
<< metal1 >>
rect -105 620 80 625
rect -105 600 -65 620
rect -45 600 80 620
rect -105 595 80 600
rect -85 230 -45 240
rect -85 210 -75 230
rect -55 210 -45 230
rect -85 200 -45 210
rect 20 230 60 240
rect 20 210 30 230
rect 50 210 60 230
rect 20 200 60 210
rect -105 -30 80 -25
rect -105 -50 -65 -30
rect -45 -50 80 -30
rect -105 -55 80 -50
<< labels >>
flabel metal1 60 -55 80 -25 1 FreeSans 200 0 0 -120 VN
port 4 n
flabel metal1 60 595 80 625 1 FreeSans 200 0 0 -120 VP
port 3 n
flabel metal1 -85 200 -45 240 1 FreeSans 200 0 0 -120 A
port 1 n
flabel metal1 20 200 60 240 1 FreeSans 200 0 0 -120 Y
port 2 n
<< end >>
