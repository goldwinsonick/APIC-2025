* PEX produced on Sun Apr 20 09:54:21 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_nand_v2.ext - technology: sky130A

.subckt goldwin_nand_v2 A B Y VP VN
X0 Y B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X2 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X3 VP B Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
C0 Y a_30_0# 0.05569f
C1 A VP 0.12847f
C2 Y VP 0.46035f
C3 a_30_0# B 0.02784f
C4 B VP 0.07186f
C5 Y A 0.0754f
C6 B A 0.15768f
C7 Y B 0.1177f
C8 Y VN 0.24822f
C9 B VN 0.37727f
C10 A VN 0.32037f
C11 VP VN 1.32377f
C12 a_30_0# VN 0.0882f
.ends

