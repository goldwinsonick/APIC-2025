* PEX produced on Sun Apr 20 09:54:22 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_mux_v2.ext - technology: sky130A

.subckt goldwin_mux_v2 A B S D VP VN
X0 goldwin_nand_v2_1.Y goldwin_not_v2_0.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X1 D goldwin_nand_v2_1.Y a_580_n370# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X2 a_580_n370# goldwin_nand_v2_3.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X3 goldwin_nand_v2_3.Y B VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X4 goldwin_not_v2_0.Y S VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X5 goldwin_not_v2_0.Y S VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X6 D goldwin_nand_v2_3.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X7 VP S goldwin_nand_v2_3.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X8 goldwin_nand_v2_3.Y S a_160_n370# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X9 goldwin_nand_v2_1.Y A a_450_130# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X10 a_160_n370# B VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X11 VP goldwin_nand_v2_1.Y D VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X12 VP A goldwin_nand_v2_1.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X13 a_450_130# goldwin_not_v2_0.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
C0 goldwin_not_v2_0.Y goldwin_nand_v2_1.Y 0.12513f
C1 D goldwin_nand_v2_1.Y 0.12616f
C2 A goldwin_nand_v2_1.Y 0.16048f
C3 D goldwin_nand_v2_3.Y 0.0895f
C4 VP goldwin_not_v2_0.Y 0.64894f
C5 VP D 0.50471f
C6 a_160_n370# S 0.03565f
C7 goldwin_nand_v2_3.Y goldwin_nand_v2_1.Y 0.20025f
C8 VP A 0.1322f
C9 A a_450_130# 0.02784f
C10 VP goldwin_nand_v2_1.Y 0.83334f
C11 a_450_130# goldwin_nand_v2_1.Y 0.07579f
C12 VP goldwin_nand_v2_3.Y 0.71027f
C13 goldwin_not_v2_0.Y S 0.16984f
C14 goldwin_nand_v2_3.Y B 0.0754f
C15 VP B 0.16956f
C16 A S 0.13502f
C17 S goldwin_nand_v2_1.Y 0.01274f
C18 a_580_n370# D 0.05569f
C19 a_160_n370# goldwin_nand_v2_3.Y 0.05569f
C20 goldwin_nand_v2_3.Y S 0.14556f
C21 a_580_n370# goldwin_nand_v2_1.Y 0.04185f
C22 VP a_160_n370# 0.01029f
C23 VP S 0.54197f
C24 A goldwin_not_v2_0.Y 0.26302f
C25 B S 0.17174f
C26 D VN 0.25653f
C27 B VN 0.34585f
C28 A VN 0.46094f
C29 S VN 1.09391f
C30 VP VN 6.18505f
C31 a_580_n370# VN 0.08205f
C32 a_160_n370# VN 0.0825f
C33 goldwin_nand_v2_3.Y VN 0.4721f
C34 a_450_130# VN 0.08821f
C35 goldwin_nand_v2_1.Y VN 0.93005f
C36 goldwin_not_v2_0.Y VN 0.49086f
.ends

