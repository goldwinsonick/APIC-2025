magic
tech sky130A
timestamp 1744280742
<< nwell >>
rect -120 175 150 515
<< nmos >>
rect -15 0 0 100
rect 50 0 65 100
<< pmos >>
rect -15 195 0 495
rect 50 195 65 495
<< ndiff >>
rect -60 85 -15 100
rect -60 15 -50 85
rect -30 15 -15 85
rect -60 0 -15 15
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 85 110 100
rect 65 15 80 85
rect 100 15 110 85
rect 65 0 110 15
<< pdiff >>
rect -60 480 -15 495
rect -60 410 -50 480
rect -30 410 -15 480
rect -60 380 -15 410
rect -60 310 -50 380
rect -30 310 -15 380
rect -60 280 -15 310
rect -60 210 -50 280
rect -30 210 -15 280
rect -60 195 -15 210
rect 0 480 50 495
rect 0 410 15 480
rect 35 410 50 480
rect 0 380 50 410
rect 0 310 15 380
rect 35 310 50 380
rect 0 280 50 310
rect 0 210 15 280
rect 35 210 50 280
rect 0 195 50 210
rect 65 480 110 495
rect 65 410 80 480
rect 100 410 110 480
rect 65 380 110 410
rect 65 310 80 380
rect 100 310 110 380
rect 65 280 110 310
rect 65 210 80 280
rect 100 210 110 280
rect 65 195 110 210
<< ndiffc >>
rect -50 15 -30 85
rect 15 15 35 85
rect 80 15 100 85
<< pdiffc >>
rect -50 410 -30 480
rect -50 310 -30 380
rect -50 210 -30 280
rect 15 410 35 480
rect 15 310 35 380
rect 15 210 35 280
rect 80 410 100 480
rect 80 310 100 380
rect 80 210 100 280
<< psubdiff >>
rect -100 85 -60 100
rect -100 15 -90 85
rect -70 15 -60 85
rect -100 0 -60 15
<< nsubdiff >>
rect -100 480 -60 495
rect -100 410 -90 480
rect -70 410 -60 480
rect -100 380 -60 410
rect -100 310 -90 380
rect -70 310 -60 380
rect -100 280 -60 310
rect -100 210 -90 280
rect -70 210 -60 280
rect -100 195 -60 210
<< psubdiffcont >>
rect -90 15 -70 85
<< nsubdiffcont >>
rect -90 410 -70 480
rect -90 310 -70 380
rect -90 210 -70 280
<< poly >>
rect -15 495 0 510
rect 50 495 65 510
rect -15 100 0 195
rect 50 100 65 195
rect -15 -65 0 0
rect 50 -65 65 0
rect -40 -75 0 -65
rect -40 -95 -30 -75
rect -10 -95 0 -75
rect -40 -105 0 -95
rect 25 -75 65 -65
rect 25 -95 35 -75
rect 55 -95 65 -75
rect 25 -105 65 -95
<< polycont >>
rect -30 -95 -10 -75
rect 35 -95 55 -75
<< locali >>
rect -100 540 -80 545
rect -100 485 -80 520
rect 90 540 110 545
rect 90 485 110 520
rect -100 480 -20 485
rect -100 410 -90 480
rect -70 410 -50 480
rect -30 410 -20 480
rect -100 380 -20 410
rect -100 310 -90 380
rect -70 310 -50 380
rect -30 310 -20 380
rect -100 280 -20 310
rect -100 210 -90 280
rect -70 210 -50 280
rect -30 210 -20 280
rect -100 205 -20 210
rect 5 480 45 485
rect 5 410 15 480
rect 35 410 45 480
rect 5 380 45 410
rect 5 310 15 380
rect 35 310 45 380
rect 5 280 45 310
rect 5 210 15 280
rect 35 210 45 280
rect 5 205 45 210
rect 70 480 110 485
rect 70 410 80 480
rect 100 410 110 480
rect 70 380 110 410
rect 70 310 80 380
rect 100 310 110 380
rect 70 280 110 310
rect 70 210 80 280
rect 100 210 110 280
rect 70 205 110 210
rect 15 150 35 205
rect 15 125 110 150
rect 90 90 110 125
rect -100 85 -20 90
rect -100 15 -90 85
rect -70 15 -50 85
rect -30 15 -20 85
rect -100 10 -20 15
rect 5 85 45 90
rect 5 15 15 85
rect 35 15 45 85
rect 5 10 45 15
rect 70 85 110 90
rect 70 15 80 85
rect 100 15 110 85
rect 70 10 110 15
rect -100 -20 -80 10
rect -100 -45 -80 -40
rect 90 -65 110 10
rect -40 -75 0 -65
rect -40 -95 -30 -75
rect -10 -95 0 -75
rect -40 -105 0 -95
rect 25 -75 65 -65
rect 25 -95 35 -75
rect 55 -95 65 -75
rect 25 -105 65 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 90 -105 130 -95
<< viali >>
rect -100 520 -80 540
rect 90 520 110 540
rect -100 -40 -80 -20
rect -30 -95 -10 -75
rect 35 -95 55 -75
rect 100 -95 120 -75
<< metal1 >>
rect -120 540 150 545
rect -120 520 -100 540
rect -80 520 90 540
rect 110 520 150 540
rect -120 515 150 520
rect -120 -20 150 -15
rect -120 -40 -100 -20
rect -80 -40 150 -20
rect -120 -45 150 -40
rect -40 -75 0 -65
rect -40 -95 -30 -75
rect -10 -95 0 -75
rect -40 -105 0 -95
rect 25 -75 65 -65
rect 25 -95 35 -75
rect 55 -95 65 -75
rect 25 -105 65 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 90 -105 130 -95
<< labels >>
flabel metal1 90 -105 130 -65 1 FreeSans 200 0 0 -120 Y
port 3 n
flabel metal1 130 -45 150 -15 1 FreeSans 200 0 0 0 VSS
port 5 n
flabel metal1 130 515 150 545 1 FreeSans 200 0 0 0 VDD
port 4 n
flabel metal1 25 -105 65 -65 1 FreeSans 200 0 0 -120 B
port 2 n
flabel metal1 -40 -105 0 -65 1 FreeSans 200 0 0 -120 A
port 1 n
<< end >>
