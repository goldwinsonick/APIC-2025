magic
tech sky130A
timestamp 1744269234
<< nwell >>
rect -110 255 735 595
<< nmos >>
rect -5 0 10 100
rect 175 0 190 100
rect 240 0 255 100
rect 375 0 390 100
rect 440 0 455 100
rect 615 0 630 100
<< pmos >>
rect -5 275 10 575
rect 175 275 190 575
rect 240 275 255 575
rect 375 275 390 575
rect 440 275 455 575
rect 615 275 630 575
<< ndiff >>
rect -50 85 -5 100
rect -50 15 -40 85
rect -20 15 -5 85
rect -50 0 -5 15
rect 10 85 55 100
rect 10 15 25 85
rect 45 15 55 85
rect 10 0 55 15
rect 130 85 175 100
rect 130 15 140 85
rect 160 15 175 85
rect 130 0 175 15
rect 190 85 240 100
rect 190 15 205 85
rect 225 15 240 85
rect 190 0 240 15
rect 255 85 300 100
rect 255 15 270 85
rect 290 15 300 85
rect 255 0 300 15
rect 330 85 375 100
rect 330 15 340 85
rect 360 15 375 85
rect 330 0 375 15
rect 390 85 440 100
rect 390 15 405 85
rect 425 15 440 85
rect 390 0 440 15
rect 455 85 500 100
rect 455 15 470 85
rect 490 15 500 85
rect 455 0 500 15
rect 570 85 615 100
rect 570 15 580 85
rect 600 15 615 85
rect 570 0 615 15
rect 630 85 675 100
rect 630 15 645 85
rect 665 15 675 85
rect 630 0 675 15
<< pdiff >>
rect -50 560 -5 575
rect -50 490 -40 560
rect -20 490 -5 560
rect -50 460 -5 490
rect -50 390 -40 460
rect -20 390 -5 460
rect -50 360 -5 390
rect -50 290 -40 360
rect -20 290 -5 360
rect -50 275 -5 290
rect 10 560 55 575
rect 10 490 25 560
rect 45 490 55 560
rect 10 460 55 490
rect 10 390 25 460
rect 45 390 55 460
rect 10 360 55 390
rect 10 290 25 360
rect 45 290 55 360
rect 10 275 55 290
rect 130 560 175 575
rect 130 490 140 560
rect 160 490 175 560
rect 130 460 175 490
rect 130 390 140 460
rect 160 390 175 460
rect 130 360 175 390
rect 130 290 140 360
rect 160 290 175 360
rect 130 275 175 290
rect 190 560 240 575
rect 190 490 205 560
rect 225 490 240 560
rect 190 460 240 490
rect 190 390 205 460
rect 225 390 240 460
rect 190 360 240 390
rect 190 290 205 360
rect 225 290 240 360
rect 190 275 240 290
rect 255 560 300 575
rect 255 490 270 560
rect 290 490 300 560
rect 255 460 300 490
rect 255 390 270 460
rect 290 390 300 460
rect 255 360 300 390
rect 255 290 270 360
rect 290 290 300 360
rect 255 275 300 290
rect 330 560 375 575
rect 330 490 340 560
rect 360 490 375 560
rect 330 460 375 490
rect 330 390 340 460
rect 360 390 375 460
rect 330 360 375 390
rect 330 290 340 360
rect 360 290 375 360
rect 330 275 375 290
rect 390 560 440 575
rect 390 490 405 560
rect 425 490 440 560
rect 390 460 440 490
rect 390 390 405 460
rect 425 390 440 460
rect 390 360 440 390
rect 390 290 405 360
rect 425 290 440 360
rect 390 275 440 290
rect 455 560 500 575
rect 455 490 470 560
rect 490 490 500 560
rect 455 460 500 490
rect 455 390 470 460
rect 490 390 500 460
rect 455 360 500 390
rect 455 290 470 360
rect 490 290 500 360
rect 455 275 500 290
rect 570 560 615 575
rect 570 490 580 560
rect 600 490 615 560
rect 570 460 615 490
rect 570 390 580 460
rect 600 390 615 460
rect 570 360 615 390
rect 570 290 580 360
rect 600 290 615 360
rect 570 275 615 290
rect 630 560 675 575
rect 630 490 645 560
rect 665 490 675 560
rect 630 460 675 490
rect 630 390 645 460
rect 665 390 675 460
rect 630 360 675 390
rect 630 290 645 360
rect 665 290 675 360
rect 630 275 675 290
<< ndiffc >>
rect -40 15 -20 85
rect 25 15 45 85
rect 140 15 160 85
rect 205 15 225 85
rect 270 15 290 85
rect 340 15 360 85
rect 405 15 425 85
rect 470 15 490 85
rect 580 15 600 85
rect 645 15 665 85
<< pdiffc >>
rect -40 490 -20 560
rect -40 390 -20 460
rect -40 290 -20 360
rect 25 490 45 560
rect 25 390 45 460
rect 25 290 45 360
rect 140 490 160 560
rect 140 390 160 460
rect 140 290 160 360
rect 205 490 225 560
rect 205 390 225 460
rect 205 290 225 360
rect 270 490 290 560
rect 270 390 290 460
rect 270 290 290 360
rect 340 490 360 560
rect 340 390 360 460
rect 340 290 360 360
rect 405 490 425 560
rect 405 390 425 460
rect 405 290 425 360
rect 470 490 490 560
rect 470 390 490 460
rect 470 290 490 360
rect 580 490 600 560
rect 580 390 600 460
rect 580 290 600 360
rect 645 490 665 560
rect 645 390 665 460
rect 645 290 665 360
<< psubdiff >>
rect -90 85 -50 100
rect -90 15 -80 85
rect -60 15 -50 85
rect -90 0 -50 15
rect 90 85 130 100
rect 90 15 100 85
rect 120 15 130 85
rect 90 0 130 15
rect 500 85 540 100
rect 500 15 510 85
rect 530 15 540 85
rect 500 0 540 15
rect 675 85 715 100
rect 675 15 685 85
rect 705 15 715 85
rect 675 0 715 15
<< nsubdiff >>
rect -90 560 -50 575
rect -90 490 -80 560
rect -60 490 -50 560
rect -90 460 -50 490
rect -90 390 -80 460
rect -60 390 -50 460
rect -90 360 -50 390
rect -90 290 -80 360
rect -60 290 -50 360
rect -90 275 -50 290
rect 90 560 130 575
rect 90 490 100 560
rect 120 490 130 560
rect 90 460 130 490
rect 90 390 100 460
rect 120 390 130 460
rect 90 360 130 390
rect 90 290 100 360
rect 120 290 130 360
rect 90 275 130 290
rect 500 560 540 575
rect 500 490 510 560
rect 530 490 540 560
rect 500 460 540 490
rect 500 390 510 460
rect 530 390 540 460
rect 500 360 540 390
rect 500 290 510 360
rect 530 290 540 360
rect 500 275 540 290
rect 675 560 715 575
rect 675 490 685 560
rect 705 490 715 560
rect 675 460 715 490
rect 675 390 685 460
rect 705 390 715 460
rect 675 360 715 390
rect 675 290 685 360
rect 705 290 715 360
rect 675 275 715 290
<< psubdiffcont >>
rect -80 15 -60 85
rect 100 15 120 85
rect 510 15 530 85
rect 685 15 705 85
<< nsubdiffcont >>
rect -80 490 -60 560
rect -80 390 -60 460
rect -80 290 -60 360
rect 100 490 120 560
rect 100 390 120 460
rect 100 290 120 360
rect 510 490 530 560
rect 510 390 530 460
rect 510 290 530 360
rect 685 490 705 560
rect 685 390 705 460
rect 685 290 705 360
<< poly >>
rect 240 620 630 635
rect -5 575 10 590
rect 175 575 190 590
rect 240 575 255 620
rect 375 575 390 590
rect 440 575 455 590
rect 615 575 630 620
rect -80 245 -40 250
rect -80 225 -70 245
rect -50 240 -40 245
rect -5 240 10 275
rect 175 250 190 275
rect 165 245 205 250
rect 165 240 175 245
rect -50 225 10 240
rect -80 220 -40 225
rect -5 100 10 225
rect 65 225 175 240
rect 195 225 205 245
rect -5 -15 10 0
rect 65 -45 80 225
rect 165 220 205 225
rect 240 195 255 275
rect 175 180 255 195
rect 175 100 190 180
rect 375 155 390 275
rect 440 160 455 275
rect 615 160 630 275
rect 215 150 390 155
rect 215 130 225 150
rect 245 140 390 150
rect 430 155 470 160
rect 245 130 255 140
rect 430 135 440 155
rect 460 135 470 155
rect 430 130 470 135
rect 615 155 660 160
rect 615 135 630 155
rect 650 135 660 155
rect 615 130 660 135
rect 215 125 255 130
rect 240 100 255 125
rect 375 100 390 115
rect 440 100 455 130
rect 615 100 630 130
rect 175 -15 190 0
rect 240 -15 255 0
rect 375 -45 390 0
rect 440 -15 455 0
rect 615 -15 630 0
rect 65 -60 390 -45
<< polycont >>
rect -70 225 -50 245
rect 175 225 195 245
rect 225 130 245 150
rect 440 135 460 155
rect 630 135 650 155
<< locali >>
rect -90 620 -70 625
rect -90 565 -70 600
rect 90 620 110 625
rect 90 565 110 600
rect 520 620 540 625
rect 520 565 540 600
rect 695 620 715 625
rect 695 565 715 600
rect -90 560 -10 565
rect -90 490 -80 560
rect -60 490 -40 560
rect -20 490 -10 560
rect -90 460 -10 490
rect -90 390 -80 460
rect -60 390 -40 460
rect -20 390 -10 460
rect -90 360 -10 390
rect -90 290 -80 360
rect -60 290 -40 360
rect -20 290 -10 360
rect -90 285 -10 290
rect 15 560 55 565
rect 15 490 25 560
rect 45 490 55 560
rect 15 460 55 490
rect 15 390 25 460
rect 45 390 55 460
rect 15 360 55 390
rect 15 290 25 360
rect 45 290 55 360
rect 15 285 55 290
rect 90 560 170 565
rect 90 490 100 560
rect 120 490 140 560
rect 160 490 170 560
rect 90 460 170 490
rect 90 390 100 460
rect 120 390 140 460
rect 160 390 170 460
rect 90 360 170 390
rect 90 290 100 360
rect 120 290 140 360
rect 160 290 170 360
rect 90 285 170 290
rect 195 560 235 565
rect 195 490 205 560
rect 225 490 235 560
rect 195 460 235 490
rect 195 390 205 460
rect 225 390 235 460
rect 195 360 235 390
rect 195 290 205 360
rect 225 290 235 360
rect 195 285 235 290
rect 260 560 300 565
rect 260 490 270 560
rect 290 490 300 560
rect 260 460 300 490
rect 260 390 270 460
rect 290 390 300 460
rect 260 360 300 390
rect 260 290 270 360
rect 290 290 300 360
rect 260 285 300 290
rect 20 250 50 285
rect -80 245 -40 250
rect -80 225 -70 245
rect -50 225 -40 245
rect -80 220 -40 225
rect 20 245 205 250
rect 20 225 175 245
rect 195 225 205 245
rect 20 220 205 225
rect 280 245 300 285
rect -75 150 -45 220
rect -75 130 -70 150
rect -50 130 -45 150
rect -75 120 -45 130
rect 20 90 50 220
rect 215 150 255 155
rect 215 130 225 150
rect 245 130 255 150
rect 215 125 255 130
rect 280 90 300 225
rect -90 85 -10 90
rect -90 15 -80 85
rect -60 15 -40 85
rect -20 15 -10 85
rect -90 10 -10 15
rect 15 85 55 90
rect 15 15 25 85
rect 45 15 55 85
rect 15 10 55 15
rect 90 85 170 90
rect 90 15 100 85
rect 120 15 140 85
rect 160 15 170 85
rect 90 10 170 15
rect 195 85 235 90
rect 195 15 205 85
rect 225 15 235 85
rect 195 10 235 15
rect 260 85 300 90
rect 260 15 270 85
rect 290 15 300 85
rect 260 10 300 15
rect 330 560 370 565
rect 330 490 340 560
rect 360 490 370 560
rect 330 460 370 490
rect 330 390 340 460
rect 360 390 370 460
rect 330 360 370 390
rect 330 290 340 360
rect 360 290 370 360
rect 330 285 370 290
rect 395 560 435 565
rect 395 490 405 560
rect 425 490 435 560
rect 395 460 435 490
rect 395 390 405 460
rect 425 390 435 460
rect 395 360 435 390
rect 395 290 405 360
rect 425 290 435 360
rect 395 285 435 290
rect 460 560 540 565
rect 460 490 470 560
rect 490 490 510 560
rect 530 490 540 560
rect 460 460 540 490
rect 460 390 470 460
rect 490 390 510 460
rect 530 390 540 460
rect 460 360 540 390
rect 460 290 470 360
rect 490 290 510 360
rect 530 290 540 360
rect 460 285 540 290
rect 570 560 610 565
rect 570 490 580 560
rect 600 490 610 560
rect 570 460 610 490
rect 570 390 580 460
rect 600 390 610 460
rect 570 360 610 390
rect 570 290 580 360
rect 600 290 610 360
rect 570 285 610 290
rect 635 560 715 565
rect 635 490 645 560
rect 665 490 685 560
rect 705 490 715 560
rect 635 460 715 490
rect 635 390 645 460
rect 665 390 685 460
rect 705 390 715 460
rect 635 360 715 390
rect 635 290 645 360
rect 665 290 685 360
rect 705 290 715 360
rect 635 285 715 290
rect 330 245 350 285
rect 330 90 350 225
rect 570 160 590 285
rect 430 155 590 160
rect 430 135 440 155
rect 460 135 590 155
rect 430 130 590 135
rect 620 155 660 160
rect 620 135 630 155
rect 650 135 660 155
rect 620 130 660 135
rect 570 90 590 130
rect 330 85 370 90
rect 330 15 340 85
rect 360 15 370 85
rect 330 10 370 15
rect 395 85 435 90
rect 395 15 405 85
rect 425 15 435 85
rect 395 10 435 15
rect 460 85 540 90
rect 460 15 470 85
rect 490 15 510 85
rect 530 15 540 85
rect 460 10 540 15
rect 570 85 610 90
rect 570 15 580 85
rect 600 15 610 85
rect 570 10 610 15
rect 635 85 715 90
rect 635 15 645 85
rect 665 15 685 85
rect 705 15 715 85
rect 635 10 715 15
rect -90 -25 -70 10
rect -90 -50 -70 -45
rect 90 -25 110 10
rect 90 -50 110 -45
rect 520 -25 540 10
rect 520 -50 540 -45
rect 695 -25 715 10
rect 695 -50 715 -45
<< viali >>
rect -90 600 -70 620
rect 90 600 110 620
rect 520 600 540 620
rect 695 600 715 620
rect 280 225 300 245
rect -70 130 -50 150
rect 225 130 245 150
rect 330 225 350 245
rect 630 135 650 155
rect -90 -45 -70 -25
rect 90 -45 110 -25
rect 520 -45 540 -25
rect 695 -45 715 -25
<< metal1 >>
rect -110 620 735 625
rect -110 600 -90 620
rect -70 600 90 620
rect 110 600 520 620
rect 540 600 695 620
rect 715 600 735 620
rect -110 595 735 600
rect 270 245 735 250
rect 270 225 280 245
rect 300 225 330 245
rect 350 225 735 245
rect 270 220 735 225
rect 620 155 735 160
rect -110 150 255 155
rect -110 130 -70 150
rect -50 130 225 150
rect 245 130 255 150
rect 620 135 630 155
rect 650 135 735 155
rect 620 130 735 135
rect -110 125 255 130
rect -110 -25 735 -20
rect -110 -45 -90 -25
rect -70 -45 90 -25
rect 110 -45 520 -25
rect 540 -45 695 -25
rect 715 -45 735 -25
rect -110 -50 735 -45
<< labels >>
rlabel metal1 -110 140 -110 140 7 A
port 1 w
rlabel metal1 735 -35 735 -35 7 VN
port 5 w
rlabel metal1 735 235 735 235 7 OUT
port 3 w
rlabel metal1 735 145 735 145 7 B
port 2 w
rlabel metal1 735 610 735 610 7 VP
port 4 w
<< end >>
