* PEX produced on Sun Apr 20 07:42:45 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from goldwin_mux_dff.ext - technology: sky130A

.subckt goldwin_mux_dff CLK A B S D Q QI VP VN
X0 goldwin_mux_0.goldwin_or_0.A a_730_650# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
X1 goldwin_mux_0.goldwin_or_0.A a_730_650# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
X2 goldwin_mux_0.goldwin_or_0.B a_1590_650# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
X3 goldwin_mux_0.goldwin_or_0.B a_1590_650# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
X4 a_730_650# A a_730_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X5 goldwin_dff_0.goldwin_nand_6.Y CLK a_3920_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X6 VP A a_730_650# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X7 VP CLK goldwin_dff_0.goldwin_nand_6.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X8 a_730_110# goldwin_mux_0.goldwin_not_0.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X9 a_3920_110# goldwin_dff_0.goldwin_not_0.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X10 a_5420_110# goldwin_dff_0.goldwin_nand_5.Y VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X11 a_730_650# goldwin_mux_0.goldwin_not_0.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X12 goldwin_dff_0.goldwin_nand_6.Y goldwin_dff_0.goldwin_not_0.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X13 Q goldwin_dff_0.goldwin_nand_5.Y VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X14 a_1590_650# B a_1590_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X15 VP B a_1590_650# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X16 a_1590_110# S VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X17 VN goldwin_mux_0.goldwin_or_0.A a_2450_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X18 a_1590_650# S VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X19 a_2450_110# goldwin_mux_0.goldwin_or_0.A a_2450_650# VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X20 Q QI a_5420_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X21 a_2450_110# goldwin_mux_0.goldwin_or_0.B VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X22 a_2450_650# goldwin_mux_0.goldwin_or_0.B VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X23 VP QI Q VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X24 D a_2450_110# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.45 ps=2.9 w=1 l=0.15
X25 a_4420_110# D VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X26 D a_2450_110# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.35 ps=6.9 w=3 l=0.15
X27 goldwin_dff_0.goldwin_nand_5.Y D VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X28 goldwin_mux_0.goldwin_not_0.Y S VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X29 goldwin_dff_0.goldwin_nand_5.Y CLK a_4420_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X30 goldwin_mux_0.goldwin_not_0.Y S VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X31 VP CLK goldwin_dff_0.goldwin_nand_5.Y VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X32 goldwin_dff_0.goldwin_not_0.Y D VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X33 QI goldwin_dff_0.goldwin_nand_6.Y a_4920_110# VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.25 ps=1.5 w=1 l=0.15
X34 goldwin_dff_0.goldwin_not_0.Y D VP VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X35 VP goldwin_dff_0.goldwin_nand_6.Y QI VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.15
X36 a_4920_110# Q VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X37 QI Q VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
C0 goldwin_mux_0.goldwin_or_0.B CLK 0.08891f
C1 goldwin_dff_0.goldwin_not_0.Y D 0.27822f
C2 CLK Q 0.02477f
C3 goldwin_mux_0.goldwin_or_0.A a_2450_650# 0.05805f
C4 CLK VP 0.21265f
C5 a_3920_110# CLK 0.03818f
C6 a_4420_110# CLK 0.02833f
C7 B CLK 0.48388f
C8 goldwin_mux_0.goldwin_or_0.B S 0.01444f
C9 a_1590_110# B 0.03383f
C10 QI a_4920_110# 0.05569f
C11 goldwin_mux_0.goldwin_not_0.Y CLK 0.0286f
C12 S VP 0.80158f
C13 a_730_110# CLK 0.02472f
C14 goldwin_dff_0.goldwin_not_0.Y CLK 0.28173f
C15 B S 0.27647f
C16 a_2450_110# D 0.11235f
C17 goldwin_mux_0.goldwin_or_0.A a_730_650# 0.10643f
C18 goldwin_mux_0.goldwin_or_0.A a_1590_650# 0.09437f
C19 goldwin_mux_0.goldwin_not_0.Y S 0.26469f
C20 goldwin_dff_0.goldwin_nand_6.Y goldwin_dff_0.goldwin_nand_5.Y 0.1456f
C21 goldwin_dff_0.goldwin_nand_6.Y QI 0.17099f
C22 goldwin_mux_0.goldwin_or_0.B a_2450_650# 0.02493f
C23 a_2450_650# VP 0.2133f
C24 a_2450_110# CLK 0.05416f
C25 A VP 0.08144f
C26 goldwin_dff_0.goldwin_nand_6.Y Q 0.20961f
C27 B A 0.24711f
C28 goldwin_dff_0.goldwin_nand_6.Y VP 0.55037f
C29 a_3920_110# goldwin_dff_0.goldwin_nand_6.Y 0.06543f
C30 a_4420_110# goldwin_dff_0.goldwin_nand_6.Y 0.03526f
C31 a_1590_650# goldwin_mux_0.goldwin_or_0.B 0.13637f
C32 goldwin_mux_0.goldwin_not_0.Y A 0.25744f
C33 a_730_110# A 0.02784f
C34 a_730_650# VP 0.54066f
C35 a_1590_650# VP 0.53929f
C36 a_730_650# B 0.06698f
C37 goldwin_dff_0.goldwin_nand_6.Y goldwin_dff_0.goldwin_not_0.Y 0.08676f
C38 a_1590_650# B 0.14514f
C39 CLK D 0.45092f
C40 goldwin_mux_0.goldwin_not_0.Y a_730_650# 0.06447f
C41 a_730_110# a_730_650# 0.05569f
C42 a_2450_110# a_2450_650# 0.19233f
C43 goldwin_mux_0.goldwin_or_0.A goldwin_mux_0.goldwin_or_0.B 0.33342f
C44 QI goldwin_dff_0.goldwin_nand_5.Y 0.37139f
C45 QI a_5420_110# 0.03661f
C46 goldwin_mux_0.goldwin_or_0.A VP 1.08145f
C47 goldwin_mux_0.goldwin_or_0.A B 0.09177f
C48 a_1590_110# CLK 0.02827f
C49 goldwin_dff_0.goldwin_nand_5.Y Q 0.51529f
C50 CLK S 0.01255f
C51 QI Q 0.48056f
C52 Q a_5420_110# 0.05569f
C53 goldwin_dff_0.goldwin_nand_5.Y VP 0.84467f
C54 QI VP 0.53693f
C55 a_4420_110# goldwin_dff_0.goldwin_nand_5.Y 0.05569f
C56 goldwin_dff_0.goldwin_nand_6.Y D 0.18595f
C57 goldwin_mux_0.goldwin_or_0.B VP 0.45811f
C58 goldwin_mux_0.goldwin_or_0.B B 0.01658f
C59 Q VP 1.17366f
C60 goldwin_mux_0.goldwin_or_0.A a_2450_110# 0.14427f
C61 B VP 0.08507f
C62 goldwin_dff_0.goldwin_nand_6.Y CLK 0.37619f
C63 goldwin_mux_0.goldwin_not_0.Y VP 0.51387f
C64 goldwin_dff_0.goldwin_not_0.Y VP 0.51422f
C65 goldwin_mux_0.goldwin_not_0.Y B 0.04556f
C66 a_730_110# B 0.03002f
C67 S A 0.16911f
C68 a_730_650# CLK 0.02849f
C69 a_1590_650# CLK 0.04269f
C70 goldwin_mux_0.goldwin_or_0.A D 0.02084f
C71 a_1590_110# a_1590_650# 0.05569f
C72 a_2450_110# goldwin_mux_0.goldwin_or_0.B 0.05068f
C73 a_730_650# S 0.09344f
C74 a_1590_650# S 0.06297f
C75 a_2450_110# VP 0.31603f
C76 goldwin_dff_0.goldwin_nand_5.Y D 0.12274f
C77 goldwin_dff_0.goldwin_nand_6.Y a_4920_110# 0.03383f
C78 goldwin_mux_0.goldwin_or_0.A CLK 0.07345f
C79 goldwin_mux_0.goldwin_or_0.A S 0.33621f
C80 CLK goldwin_dff_0.goldwin_nand_5.Y 0.12095f
C81 a_730_650# A 0.13804f
C82 D VP 1.08609f
C83 QI VN 0.77397f
C84 Q VN 0.65094f
C85 CLK VN 3.17317f
C86 D VN 1.0138f
C87 B VN 0.72065f
C88 A VN 0.40106f
C89 S VN 0.87238f
C90 VP VN 13.6975f
C91 a_5420_110# VN 0.08711f
C92 a_4920_110# VN 0.08755f
C93 a_4420_110# VN 0.08572f
C94 a_3920_110# VN 0.08755f
C95 a_1590_110# VN 0.07692f
C96 a_730_110# VN 0.07692f
C97 a_2450_650# VN 0.01525f
C98 goldwin_dff_0.goldwin_nand_5.Y VN 0.58442f
C99 goldwin_dff_0.goldwin_nand_6.Y VN 0.93533f
C100 goldwin_dff_0.goldwin_not_0.Y VN 0.54656f
C101 a_2450_110# VN 0.64876f
C102 goldwin_mux_0.goldwin_or_0.A VN 0.59629f
C103 goldwin_mux_0.goldwin_or_0.B VN 0.64107f
C104 a_1590_650# VN 0.55852f
C105 a_730_650# VN 0.55835f
C106 goldwin_mux_0.goldwin_not_0.Y VN 0.55349f
.ends

