magic
tech sky130A
timestamp 1744387960
<< nwell >>
rect -105 250 145 590
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
<< pmos >>
rect 0 270 15 570
rect 65 270 80 570
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 125 100
rect 80 15 95 85
rect 115 15 125 85
rect 80 0 125 15
<< pdiff >>
rect -45 555 0 570
rect -45 485 -35 555
rect -15 485 0 555
rect -45 455 0 485
rect -45 385 -35 455
rect -15 385 0 455
rect -45 355 0 385
rect -45 285 -35 355
rect -15 285 0 355
rect -45 270 0 285
rect 15 555 65 570
rect 15 485 30 555
rect 50 485 65 555
rect 15 455 65 485
rect 15 385 30 455
rect 50 385 65 455
rect 15 355 65 385
rect 15 285 30 355
rect 50 285 65 355
rect 15 270 65 285
rect 80 555 125 570
rect 80 485 95 555
rect 115 485 125 555
rect 80 455 125 485
rect 80 385 95 455
rect 115 385 125 455
rect 80 355 125 385
rect 80 285 95 355
rect 115 285 125 355
rect 80 270 125 285
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
<< pdiffc >>
rect -35 485 -15 555
rect -35 385 -15 455
rect -35 285 -15 355
rect 30 485 50 555
rect 30 385 50 455
rect 30 285 50 355
rect 95 485 115 555
rect 95 385 115 455
rect 95 285 115 355
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
<< nsubdiff >>
rect -85 555 -45 570
rect -85 485 -75 555
rect -55 485 -45 555
rect -85 455 -45 485
rect -85 385 -75 455
rect -55 385 -45 455
rect -85 355 -45 385
rect -85 285 -75 355
rect -55 285 -45 355
rect -85 270 -45 285
<< psubdiffcont >>
rect -75 15 -55 85
<< nsubdiffcont >>
rect -75 485 -55 555
rect -75 385 -55 455
rect -75 285 -55 355
<< poly >>
rect 0 570 15 585
rect 65 570 80 585
rect -85 220 -45 225
rect 0 220 15 270
rect -85 200 -75 220
rect -55 200 15 220
rect -85 195 -45 200
rect 0 100 15 200
rect 65 160 80 270
rect 40 155 80 160
rect 40 135 50 155
rect 70 135 80 155
rect 40 130 80 135
rect 65 100 80 130
rect 0 -15 15 0
rect 65 -15 80 0
<< polycont >>
rect -75 200 -55 220
rect 50 135 70 155
<< locali >>
rect -65 620 -45 625
rect -65 560 -45 600
rect 85 620 105 625
rect 85 560 105 600
rect -85 555 -5 560
rect -85 485 -75 555
rect -55 485 -35 555
rect -15 485 -5 555
rect -85 455 -5 485
rect -85 385 -75 455
rect -55 385 -35 455
rect -15 385 -5 455
rect -85 355 -5 385
rect -85 285 -75 355
rect -55 285 -35 355
rect -15 285 -5 355
rect -85 280 -5 285
rect 20 555 60 560
rect 20 485 30 555
rect 50 485 60 555
rect 20 455 60 485
rect 20 385 30 455
rect 50 385 60 455
rect 20 355 60 385
rect 20 285 30 355
rect 50 285 60 355
rect 20 280 60 285
rect 85 555 125 560
rect 85 485 95 555
rect 115 485 125 555
rect 85 455 125 485
rect 85 385 95 455
rect 115 385 125 455
rect 85 355 125 385
rect 85 285 95 355
rect 115 285 125 355
rect 85 280 125 285
rect -85 220 -45 230
rect -85 200 -75 220
rect -55 200 -45 220
rect 30 220 50 280
rect 85 220 125 230
rect 30 200 95 220
rect 115 200 125 220
rect -85 190 -45 200
rect 85 190 125 200
rect -85 155 -45 165
rect 40 155 80 160
rect -85 135 -75 155
rect -55 135 50 155
rect 70 135 80 155
rect -85 125 -45 135
rect 40 130 80 135
rect 105 90 125 190
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect 85 85 125 90
rect 85 15 95 85
rect 115 15 125 85
rect 85 10 125 15
rect -65 -30 -45 10
rect -65 -55 -45 -50
<< viali >>
rect -65 600 -45 620
rect 85 600 105 620
rect -75 200 -55 220
rect 95 200 115 220
rect -75 135 -55 155
rect -65 -50 -45 -30
<< metal1 >>
rect -105 620 145 625
rect -105 600 -65 620
rect -45 600 85 620
rect 105 600 145 620
rect -105 595 145 600
rect -85 220 -45 230
rect -85 200 -75 220
rect -55 200 -45 220
rect -85 190 -45 200
rect 85 220 125 230
rect 85 200 95 220
rect 115 200 125 220
rect 85 190 125 200
rect -85 155 -45 165
rect -85 135 -75 155
rect -55 135 -45 155
rect -85 125 -45 135
rect -105 -30 145 -25
rect -105 -50 -65 -30
rect -45 -50 145 -30
rect -105 -55 145 -50
<< labels >>
flabel metal1 -85 190 -45 230 1 FreeSans 200 0 0 -120 A
port 1 n
flabel metal1 -85 125 -45 165 1 FreeSans 200 0 0 -120 B
port 2 n
flabel metal1 85 190 125 230 1 FreeSans 200 0 0 -120 Y
port 3 n
flabel metal1 125 595 145 625 1 FreeSans 200 0 0 -120 VP
port 4 n
flabel metal1 125 -55 145 -25 1 FreeSans 200 0 0 -120 VN
port 5 n
<< end >>
